module router_sync(
	input clk,resetn,detect_add,full_0,full_1,full_2,empty_0,empty_1,empty_2,write_enb_reg,read_enb_0,read_enb_1,read_enb_2,
	input [1:0] data_in,
	output reg  [2:0]write_enb,
	output reg fifo_full,soft_reset_0,soft_reset_1,soft_reset_2,
	output vld_out_0,vld_out_1,vld_out_2
	);
	
	reg [1:0]addr;
	reg [4:0] count_0,count_1,count_2;
	
	//write_enb block
  always@(posedge clk)
		if(!resetn)
			addr<=2'b00;
		else if(detect_add==1)
			addr<=data_in;
		else
			addr<=addr;
			
  always@(addr,write_enb_reg )
		if(write_enb_reg==1)
			case(addr)
				2'b00: write_enb=3'b001;
				2'b01: write_enb=3'b010;
				2'b10: write_enb=3'b100;
				default : write_enb=3'b000;
			endcase
		else 
			write_enb=3'b000;
			
	//fifo full block
	always@(*)
		case(addr)
				2'b00: fifo_full=full_0?1:0;
				2'b01: fifo_full=full_1?1:0;
				2'b10: fifo_full=full_2?1:0;
				default : fifo_full=0;
		endcase
	
	//count for soft_rest_signal
	always@(posedge clk)
		if(!resetn)
			begin
			count_0<=1;
			soft_reset_0<=0;
			end
		else if(vld_out_0==0)
			count_0<=1;
		else if(read_enb_0==1)
			count_0<=1;
		else if(count_0==30)
			begin
			count_0<=1;
			soft_reset_0<=1;
			end
		else
			begin
			count_0<=count_0+1;
			soft_reset_0<=0;
			end

	always@(posedge clk)
		if(!resetn)
			begin
			count_1<=1;
			soft_reset_1<=0;
			end
		else if(vld_out_1==0)
			count_1<=1;
		else if(read_enb_1==1)
			count_1<=1;
		else if(count_1==30)
			begin
			count_1<=1;
			soft_reset_1<=1;
			end
		else
			begin
			count_1<=count_1+1;
			soft_reset_1<=0;
			end

	always@(posedge clk)
		if(!resetn)
			begin
			count_2<=1;
			soft_reset_2<=0;
			end
		else if(vld_out_2==0)
			count_2<=1;
		else if(read_enb_2==1)
			count_2<=1;
		else if(count_2==30)
			begin
			count_2<=1;
			soft_reset_2<=1;
			end
		else
			begin
			count_2<=count_2+1;
			soft_reset_2<=0;
			end


	//vld_out signal
	assign vld_out_0=~empty_0;
	assign vld_out_1=~empty_1;
	assign vld_out_2=~empty_2;
	
endmodule
